module top_v1
  #(parameter random = 16,
  parameter blah = 2)
  (
   input CLK, 
   input RST,
   input toot,
   input enable,
   input [random:0] value,
   output [7:0] led
  );
  reg [31:0] count;
  reg [7:0] state;
  assign led = count[23:16];
  always @(posedge CLK) begin
    if(RST) begin
      count <= 0;
      state <= 0;
    end else begin
      if(state == 0) begin
        if(enable) state <= 1;
      end else if(state == 1) begin
        state <= 2;
      end else if(state == 2) begin
        count <= count + value;
        state <= 0;
      end
    end
  end
  blink inst_1 (.CLK(CLK));
  test inst_2 ();
  moduleName inst_3 ();

endmodule
