module static (
    input something
);
    
endmodule
